module pll (
  input                   refclk,
  input                   rst,
  output                  outclk_0 /* verilator public */, 
  output                  outclk_1  /* verilator public */, 
  output                  locked
);

endmodule
