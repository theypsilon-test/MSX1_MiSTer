// WD279x FDC
//
// Copyright (c) 2024-2025 Molekula
//
// All rights reserved
//
// Redistribution and use in source and synthezised forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// * Redistributions of source code must retain the above copyright notice,
//   this list of conditions and the following disclaimer.
//
// * Redistributions in synthesized form must reproduce the above copyright
//   notice, this list of conditions and the following disclaimer in the
//   documentation and/or other materials provided with the distribution.
//
// * Neither the name of the author nor the names of other contributors may
//   be used to endorse or promote products derived from this software without
//   specific prior written agreement from the author.
//
// * License is granted for non-commercial use only.  A fee may not be charged
//   for redistributions as source code or in synthesized/hardware form without
//   specific prior written agreement from the author.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
// THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR
// PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE AUTHOR OR CONTRIBUTORS BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
// INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
// CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.
//

module wd279x_command_IV 
(
	input  logic        clk,         // sys clock
	output logic        interrupt,
	input  logic        MRn,	     // master reset
	input  logic        command_start,
	input  logic  [7:0] command,
	output logic  [7:0] status,
	output logic        INTRQ,
	input  logic        INTRQ_ACK,
	input  logic 		INDEXn,
	input  logic        READYn,
	input  logic 		WPROTn,
	input  logic 		TRK00n,
	input  logic        HLD
);

	assign status = command[7:4] != 4'hD ? 8'h00 : {READYn, ~WPROTn, HLD, 1'b0, 1'b0, ~TRK00n, ~INDEXn, 1'b0};

	logic last_READY;
	always_ff @(posedge clk) begin
		last_READY <= READYn;
		interrupt <= 0;
		
		if (~MRn) begin
			INTRQ <= 0;
		end else begin
			if (command_start) INTRQ <= 0;

			if (INTRQ_ACK) INTRQ <= 0;

			if (command[7:4] == 4'hD) begin
				if (command_start) begin
					$display("Command IV Command %x %t", command, $time);
					INTRQ <= command[3];
					interrupt <= 1;
				end
				if (command[0] && !READYn && last_READY) INTRQ <= 1;
				if (command[1] && READYn && !last_READY) INTRQ <= 1;
				if (command[2] && !INDEXn) INTRQ <= 1;
			end
		end
	end
endmodule

