/*verilator tracing_off*/
module opll
(
   input clk,
   input cen,
   input rst,
   input [7:0] din,
   input addr,
   input [2:0] wr,
   input [2:0] cs,
   output signed [15:0] sound
);


endmodule