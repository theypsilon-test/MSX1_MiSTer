   module msx #(parameter sysCLK)
(
   input                    core_reset,
   input                    core_hard_reset,
   //Clock
   clock_bus_if.base_mp     clock_bus,
   //Video
   video_bus_if.device_mp   video_bus,
   vram_bus_if.device_mp    vram_bus,
   //Ext SD card
   ext_sd_card_if.device_mp ext_SD_card_bus,
   //Flash acces to SDRAM
   flash_bus_if.device_mp   flash_bus,
   //debug
   output MSX::cpu_regs_t   cpu_regs,
   output  [31:0]           opcode,
   output  [1:0]            opcode_num,
   output                   opcode_out,
   output logic [15:0]      opcode_PC_start,
   //I/O
   output            [15:0] audio_L,
   output            [15:0] audio_R,
   input             [10:0] ps2_key,
   input              [5:0] joy[2],
   //Cassete
   output                   tape_motor_on,
   input                    tape_in,
   //MSX config
   input             [64:0] rtc_time,
   input MSX::user_config_t msx_user_config,
   input                    sram_save,
   input                    sram_load,
   //IOCTL
   input                    ioctl_download,
   input             [15:0] ioctl_index,
   input             [26:0] ioctl_addr,
   //SDRAM/BRAM
   output            [26:0] ram_addr,
   output             [7:0] ram_din,
   output                   ram_rnw,
   output                   sdram_ce,
   output                   bram_ce,
   input              [7:0] ram_dout,
   input              [1:0] sdram_size,
   input MSX::slot_expander_t slot_expander[4],
   input MSX::block_t       slot_layout[64],
   input MSX::lookup_RAM_t  lookup_RAM[16],
   input MSX::lookup_SRAM_t lookup_SRAM[4],
   input MSX::io_device_t   io_device[32][3],
   input MSX::io_device_mem_ref_t io_memory[8],
   input MSX::msx_config_t  msx_config,
   //KBD
   input MSX::kb_memory_t   kb_upload_memory,
   //SD FDC
   FDD_if.FDC_mp           FDD_bus[3],
   
   /*
   input                    img_mounted,
   input             [31:0] img_size,
   input                    img_readonly,
   output            [31:0] sd_lba,
   output                   sd_rd,
   output                   sd_wr,
   input                    sd_ack,
   input             [13:0] sd_buff_addr,
   input              [7:0] sd_buff_dout,
   output             [7:0] sd_buff_din,
   input                    sd_buff_wr
);

device_bus device_bus();
cpu_bus_if cpu_bus(clock_bus.clk, reset);

//  -----------------------------------------------------------------------------
//  -- reset
//  -----------------------------------------------------------------------------
   logic reset = '0;
   always_ff @(posedge clock_bus.clk) begin
      reset <= core_hard_reset || (core_reset && ~reset_lock) || reset_request;
   end

//  -----------------------------------------------------------------------------
//  -- Audio MIX
//  -----------------------------------------------------------------------------
wire [15:0] compr_L[7:0], compr_R[7:0];
wire  [9:0] sysAudio    = {4'b0, keybeep,5'b00000} + {5'b0, (tape_in & ~tape_motor_on),4'b0000};
wire [16:0] fm          = {3'b00, sysAudio, 4'b0000};
wire [16:0] audio_mix_L   = {device_sound_L[15], device_sound_L} + fm;
wire [16:0] audio_mix_R   = {device_sound_R[15], device_sound_R} + fm;
assign compr_L            = '{ {1'b1, audio_mix_L[13:0], 1'b0}, 16'h8000, 16'h8000, 16'h8000, 16'h7FFF, 16'h7FFF, 16'h7FFF,  {1'b0, audio_mix_L[13:0], 1'b0}};
assign compr_R            = '{ {1'b1, audio_mix_R[13:0], 1'b0}, 16'h8000, 16'h8000, 16'h8000, 16'h7FFF, 16'h7FFF, 16'h7FFF,  {1'b0, audio_mix_R[13:0], 1'b0}};
assign audio_L            = compr_L[audio_mix_L[16:14]];
assign audio_R            = compr_R[audio_mix_R[16:14]];

//  -----------------------------------------------------------------------------
//  -- T80 CPU
//  -----------------------------------------------------------------------------
wire [7:0] d_to_cpu;
wire cpu_interrupt;


logic cpu_clk;
always_comb begin
   case(cpu_clock_sel)
      2'b00: cpu_clk = clock_bus.ce_3m58_n;
      2'b01: cpu_clk = clock_bus.ce_10m7_n;
      2'b10: cpu_clk = clock_bus.ce_5m39_n;
      2'b11: cpu_clk = clock_bus.ce_3m58_n;
      endcase
end
wire m1_n, mreq_n, iorq_n, rd_n, wr_n, rfsh_n;

assign cpu_bus.cpu_mp.mreq    = ~mreq_n;
assign cpu_bus.cpu_mp.iorq    = ~iorq_n;
assign cpu_bus.cpu_mp.m1      = ~m1_n;
assign cpu_bus.cpu_mp.rd      = ~rd_n;
assign cpu_bus.cpu_mp.wr      = ~wr_n;
assign cpu_bus.cpu_mp.rfsh    = ~rfsh_n;
assign cpu_bus.cpu_mp.cpu_clk = cpu_clk;
assign cpu_bus.cpu_mp.req     = ~((iorq_n & mreq_n) | (wr_n & rd_n) | iack);

logic iack;
always @(posedge cpu_bus.clk) begin
   if (cpu_bus.reset) 
   iack <= 0;
   else begin
   if (iorq_n && mreq_n)
      iack <= 0;
   else
      if (cpu_bus.cpu_mp.req)
         iack <= 1;
   end
end
  

TV80a #(.Mode(0), .R800_MULU(1), .IOWait(1)) Z80
(
   .RESET_n(~reset),
   .R800_mode('0),
   .CLK_n(cpu_clk),
   .WAIT_n(wait_n),
   .INT_n(~cpu_interrupt),
   .NMI_n('1),
   .BUSRQ_n('1),
   .M1_n(m1_n),
   .MREQ_n(mreq_n),
   .IORQ_n(iorq_n),
   .RD_n(rd_n),
   .WR_n(wr_n),
   .RFSH_n(rfsh_n),
   .HALT_n(),
   .BUSAK_n(),
   .A(cpu_bus.cpu_mp.addr),
   .DI(d_to_cpu),
   .DO(cpu_bus.cpu_mp.data)
);
//  -----------------------------------------------------------------------------
//  -- WAIT CPU
//  -----------------------------------------------------------------------------
logic wait_n, dev_cpu_wait;
logic [2:0] wait_count = 0;
logic last_m1;

always_ff @(negedge cpu_bus.cpu_clk) begin
   last_m1 <= cpu_bus.device_mp.m1;
   if (~last_m1 && cpu_bus.device_mp.m1) begin
      wait_count <= msx_config.wait_count;
   end else if (wait_count != 3'd0) begin
      wait_count <= wait_count - 3'b01;
   end
end

assign wait_n = wait_count == 3'd00 && ~dev_cpu_wait;

//  -----------------------------------------------------------------------------
//  -- Slots 
//  -----------------------------------------------------------------------------
wire [1:0] active_slot;

assign active_slot =    //~map_valid                             ? default_slot   :
                        cpu_bus.device_mp.addr[15:14] == 2'b00 ? slot_config[1:0] :
                        cpu_bus.device_mp.addr[15:14] == 2'b01 ? slot_config[3:2] :
                        cpu_bus.device_mp.addr[15:14] == 2'b10 ? slot_config[5:4] :
                                                                 slot_config[7:6] ;

//  -----------------------------------------------------------------------------
//  -- CPU data multiplex
//  -----------------------------------------------------------------------------
assign d_to_cpu = ~cpu_bus.device_mp.rd   ? 8'hFF           :
                  device_oe_rq            ? device_data     :                       // Prioritní data.
                  slot_oe_rq              ? d_from_slots    :                       // Prioritní data.
                                            device_data & ram_dout & d_from_slots;

wire signed [15:0] device_sound_L, device_sound_R;

assign ram_addr = slots_ram_addr & device_ram_addr;
assign sdram_ce = slots_ram_ce   | device_ram_ce;

wire  [7:0] device_data;
wire  [7:0] data_to_mapper;
wire  [7:0] slot_config;
wire [26:0] device_ram_addr;
wire        device_ram_ce;
wire        device_oe_rq;
wire        keybeep;
wire        reset_lock, reset_request, ocm_megaSD_enable;
wire [1:0]  ocm_slot2_mode;
wire        ocm_slot1_mode;
wire [1:0]  cpu_clock_sel;
devices #(.sysCLK(sysCLK)) devices
(
   .clock_bus(clock_bus),
   .cpu_bus(cpu_bus),
   .device_bus(device_bus),
   .FDD_bus(FDD_bus),
   .io_device(io_device),
   .io_memory(io_memory),
   .sound_L(device_sound_L),
   .sound_R(device_sound_R),
   .data(device_data),
   .data_oe_rq(device_oe_rq),
   .data_to_mapper(data_to_mapper),
   .ram_cs(device_ram_ce),
   .ram_addr(device_ram_addr),
   .vram_bus(vram_bus),
   .video_bus(video_bus),
   .cpu_interrupt(cpu_interrupt),
   .kb_upload_memory(kb_upload_memory),
   .ps2_key(ps2_key),
   .rtc_time(rtc_time),
   .joy(joy),
   .tape_in(tape_in),
   .tape_motor_on(tape_motor_on),
   .slot_config(slot_config),
   .keybeep(keybeep),
   .msx_user_config(msx_user_config),
   .reset_lock(reset_lock),
   .reset_request(reset_request),
   .cpu_wait(dev_cpu_wait),
   .cpu_clock_sel(cpu_clock_sel),
   .ocm_megaSD_enable(ocm_megaSD_enable),
   .ocm_slot1_mode(ocm_slot1_mode),
   .ocm_slot2_mode(ocm_slot2_mode)
);

wire  [7:0] d_from_slots;
wire [26:0] slots_ram_addr;
wire        slots_ram_ce;
wire        slot_oe_rq;
msx_slots msx_slots
(
   .clock_bus(clock_bus),
   .cpu_bus(cpu_bus),
   .device_bus(device_bus),
   .ext_SD_card_bus(ext_SD_card_bus),
   .flash_bus(flash_bus),
   .slot_expander(slot_expander),
   .slot_layout(slot_layout),
   .lookup_RAM(lookup_RAM),
   .lookup_SRAM(lookup_SRAM),
   .data(d_from_slots),
   .data_oe_rq(slot_oe_rq),
   .ram_addr(slots_ram_addr),
   .ram_din(ram_din),
   .ram_rnw(ram_rnw),
   .ram_dout(ram_dout),
   .sdram_ce(slots_ram_ce),
   .bram_ce(bram_ce),
   .sdram_size(sdram_size),
   .active_slot(active_slot),
   .data_to_mapper(data_to_mapper),
   .ocm_megaSD_enable(ocm_megaSD_enable),
   .ocm_slot1_mode(ocm_slot1_mode),
   .ocm_slot2_mode(ocm_slot2_mode)
);

endmodule
