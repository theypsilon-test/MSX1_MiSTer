/*verilator tracing_off*/
module mapper_gamemaster2 (
    cpu_bus     cpu_bus,   // Interface for CPU communication
    mapper_out  out,       // Interface for mapper output
    mapper      mapper     // Struct containing mapper configuration and parameters
);

    // Memory mapping control signals
    wire cs, mapper_en, rom_mapped;

    // Enable mapper if the mapper type is GameMaster2
    assign mapper_en = (mapper.typ == MAPPER_GM2);

    // Determine if the ROM is mapped (address range 4000h - BFFFh)
    assign rom_mapped = cpu_bus.addr[15] ^ cpu_bus.addr[14];

    // Chip select (cs) is active if the mapper is enabled and the CPU is performing a memory request (mreq)
    assign cs = mapper_en && cpu_bus.mreq;

    // Bank registers for memory mapping
    logic [5:0] bank1, bank2, bank3;

    // Bank switching logic based on CPU reset and clock signals
    always @(posedge cpu_bus.reset or posedge cpu_bus.clk) begin
        if (cpu_bus.reset) begin
            // Initialize banks after reset
            bank1 <= 6'h01;  // Default bank 1
            bank2 <= 6'h02;  // Default bank 2
            bank3 <= 6'h03;  // Default bank 3
        end else begin
            if (cs && cpu_bus.wr) begin
                // Update bank registers based on the address range during a write
                case (cpu_bus.addr[15:12])
                    4'h6: bank1 <= cpu_bus.data[5:0];  // Bank 1 (6000h - 6FFFh)
                    4'h8: bank2 <= cpu_bus.data[5:0];  // Bank 2 (8000h - 8FFFh)
                    4'hA: bank3 <= cpu_bus.data[5:0];  // Bank 3 (A000h - AFFFh)
                    default: ;  // No action for other address ranges
                endcase
            end
        end
    end

    // Bank selection logic based on the CPU address range
    wire [5:0] bank_base = (cpu_bus.addr[15:13] == 3'b010) ? 6'h00 :  // Fixed bank for 4000h - 5FFFh
                           (cpu_bus.addr[15:13] == 3'b011) ? bank1 :  // Bank 1 (6000h - 7FFFh)
                           (cpu_bus.addr[15:13] == 3'b100) ? bank2 :  // Bank 2 (8000h - 9FFFh)
                                                             bank3 ;  // Bank 3 (A000h - BFFFh)

    // Generate RAM and SRAM addresses based on the selected bank and CPU address
    wire [26:0] ram_addr  = {10'b0, bank_base[3:0], cpu_bus.addr[12:0]};  // RAM address
    wire [26:0] sram_addr = {14'b0, bank_base[5],   cpu_bus.addr[11:0]};  // SRAM address

    // Enable SRAM if bit 4 of the bank register is set; otherwise, enable RAM for read operations
    wire sram_en = bank_base[4];
    wire ram_en  = ~sram_en && cpu_bus.rd && rom_mapped;

    // Output control signals
    assign out.sram_cs = cs && sram_en;  // SRAM chip select
    assign out.ram_cs  = cs && ram_en;   // RAM chip select
    assign out.rnw     = ~(out.sram_cs && cpu_bus.wr && cpu_bus.addr[15:12] == 4'hB);  // Read/Write control signal
    assign out.addr    = cs ? (sram_en ? sram_addr : ram_addr) : {27{1'b1}};  // Address output, default to all 1s if not selected

endmodule
