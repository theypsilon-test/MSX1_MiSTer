module top
(
   input sclk              /* verilator public */,
   input fclk              /* verilator public */,
   input rstn              /* verilator public */,
   input RDn               /* verilator public */,
   input WRn               /* verilator public */,
   input CSn               /* verilator public */,
   input A0                /* verilator public */,
   input [7:0] WDAT        /* verilator public */,
   output [7:0] RDAT       /* verilator public */,
   output DATOE            /* verilator public */,
   input DACKn             /* verilator public */,
   output DRQ              /* verilator public */,
   input  TC               /* verilator public */,
   output INTn             /* verilator public */,
   input WAITIN            /* verilator public */,

   // Mister IMAGE
   input   [5:0] img_mounted    /* verilator public */,
   input  [63:0] img_size       /* verilator public */,

   //SD block level access
   output logic [31:0] sd_lba[6]      /* verilator public */,
   output  [5:0] sd_blk_cnt[6]  /* verilator public */,
   output  logic [5:0] sd_rd          /* verilator public */,
   output  [5:0] sd_wr          /* verilator public */,
   input   [5:0] sd_ack         /* verilator public */,
   
   // SD byte level access. Signals for 2-PORT altsyncram.
   input  [13:0] sd_buff_addr   /* verilator public */,
   input   [7:0] sd_buff_dout   /* verilator public */,
   output  [7:0] sd_buff_din[6] /* verilator public */,
   input         sd_buff_wr     /* verilator public */
);

initial begin
   sd_lba = '{32'd0, 32'd0, 32'd0, 32'd0, 32'd0, 32'd0};
   sd_rd = 6'b0;
end

logic [3:0] cnt = 4'd1;
logic last_mount = 0;
always_ff @(posedge fclk) begin
   if (!last_mount && img_mounted[3]) begin
      cnt <= '1;
   end else begin
      if (img_mounted[3]) begin
         if (cnt > '0) begin
            cnt <= cnt - 1'b1;
         end else begin
            sd_lba[3] <= 32'd1;
            sd_rd[3] <= '1;
         end
      end
   end
   last_mount <= img_mounted[3];
end

tc8566af tc8566af (
   .RDn(RDn),
   .WRn(WRn),
   .CSn(CSn),
   .A0(A0),
   .WDAT(WDAT),
   .RDAT(RDAT),
   .DATOE(DATOE),
   .DACKn(DACKn),
   .DRQ(DRQ),
   .TC(TC),
   .INTn(INTn),
   .WAITIN(WAITIN),

   .WREN(),
   .WRBIT(),
   .RDBIT(),
   .STEP(),
   .SDIR(),
   .WPRT(),
   .track0(),
   .index(),
   .side(),
   .usel(),
   .READY(),
   .TWOSIDE(),

   .int0(),
   .int1(),
   .int2(),
   .int3(),

   .td0(),
   .td1(),
   .td2(),
   .td3(),

   .hmssft(),
   
   .busy(),
   .mfm(),

   .ismode(),

   .sclk(sclk),
   .fclk(fclk),
   .rstn(rstn)
);

endmodule