/*verilator tracing_off*/
module devices (
    cpu_bus         cpu_bus,            // Interface for CPU communication
    device_bus      device_bus,         // Interface for device control
    input     [2:0] dev_enable[0:(1 << $bits(device_t))-1], // Enable signals for each device
    input MSX::io_device_t   io_device[16],  // Array of IO devices with port and mask info
    input     [7:0] dev_dout,           // Data output from device
    input           dev_rd,             // Read request signal
    output signed [15:0] sound          // Combined sound output
);

    // Combine sound outputs from the enabled OPL3 channels
    assign sound = (dev_enable[DEV_OPL3][0] ? sound_OPL3[0] : '0) +
                   (dev_enable[DEV_OPL3][1] ? sound_OPL3[1] : '0) +
                   (dev_enable[DEV_OPL3][2] ? sound_OPL3[2] : '0);

    // IO operation signal
    wire io_op = cpu_bus.iorq && ~cpu_bus.m1;

    // Enable signals for OPL3
    wire [2:0] opl3_en; 
    io_decoder #(.DEV_NAME(DEV_OPL3)) opl_decoder (
        .cpu_addr(cpu_bus.addr[7:0]),
        .io_device(io_device),
        .enable(opl3_en)
    );

    // OPL3 instances for sound generation
    wire signed [15:0] sound_OPL3[0:2];
    logic [2:0] opl3_enabled;
    genvar i;

    generate
        for (i = 0; i < 3; i++) begin : OPL3_INSTANCES
            jt2413 OPL3_i (
                .clk(cpu_bus.clk),
                .rst(cpu_bus.reset),
                .cen(cpu_bus.clk_en),
                .din(cpu_bus.data),
                .addr(cpu_bus.addr[0]),
                .cs_n(~(io_op && opl3_en[i] && opl3_enabled[i])),  // Chip select for OPL3
                .wr_n(~(cpu_bus.wr | device_bus.we)),              // Write enable
                .snd(sound_OPL3[i]),                               // Sound output
                .sample()                                          // Sample output (unused)
            );
        end
    endgenerate

    // Control logic for enabling or disabling OPL3 channels
    always @(posedge cpu_bus.clk) begin
        if (cpu_bus.reset) begin
            // Default to all OPL3 channels enabled
            opl3_enabled <= 3'b111;
        end else if (device_bus.typ == DEV_OPL3 && device_bus.num < 3) begin
            // Update enabled status for the specific OPL3 channel
            opl3_enabled[device_bus.num] <= device_bus.en;
        end
    end

endmodule

module io_decoder (
    input  logic [7:0]           cpu_addr,     // Address from CPU bus
    input  MSX::io_device_t      io_device[16],// Array of IO devices
    output logic [2:0]           enable        // Enable signals for devices
);
    parameter DEV_NAME;

    // Generate enable signal based on matching CPU address and IO device information
    assign enable = 
                      ((cpu_addr & io_device[0].mask) == io_device[0].port && io_device[0].id == DEV_NAME ? (3'b001 << io_device[0].num) : 3'b000) |
                      ((cpu_addr & io_device[1].mask) == io_device[1].port && io_device[1].id == DEV_NAME ? (3'b001 << io_device[1].num) : 3'b000) |
                      ((cpu_addr & io_device[2].mask) == io_device[2].port && io_device[2].id == DEV_NAME ? (3'b001 << io_device[2].num) : 3'b000) |
                      ((cpu_addr & io_device[3].mask) == io_device[3].port && io_device[3].id == DEV_NAME ? (3'b001 << io_device[3].num) : 3'b000) |
                      ((cpu_addr & io_device[4].mask) == io_device[4].port && io_device[4].id == DEV_NAME ? (3'b001 << io_device[4].num) : 3'b000) |
                      ((cpu_addr & io_device[5].mask) == io_device[5].port && io_device[5].id == DEV_NAME ? (3'b001 << io_device[5].num) : 3'b000) |
                      ((cpu_addr & io_device[6].mask) == io_device[6].port && io_device[6].id == DEV_NAME ? (3'b001 << io_device[6].num) : 3'b000) |
                      ((cpu_addr & io_device[7].mask) == io_device[7].port && io_device[7].id == DEV_NAME ? (3'b001 << io_device[7].num) : 3'b000) |
                      ((cpu_addr & io_device[8].mask) == io_device[8].port && io_device[8].id == DEV_NAME ? (3'b001 << io_device[8].num) : 3'b000) |
                      ((cpu_addr & io_device[9].mask) == io_device[9].port && io_device[9].id == DEV_NAME ? (3'b001 << io_device[9].num) : 3'b000) |
                      ((cpu_addr & io_device[10].mask) == io_device[10].port && io_device[10].id == DEV_NAME ? (3'b001 << io_device[10].num) : 3'b000) |
                      ((cpu_addr & io_device[11].mask) == io_device[11].port && io_device[11].id == DEV_NAME ? (3'b001 << io_device[11].num) : 3'b000) |
                      ((cpu_addr & io_device[12].mask) == io_device[12].port && io_device[12].id == DEV_NAME ? (3'b001 << io_device[12].num) : 3'b000) |
                      ((cpu_addr & io_device[13].mask) == io_device[13].port && io_device[13].id == DEV_NAME ? (3'b001 << io_device[13].num) : 3'b000) |
                      ((cpu_addr & io_device[14].mask) == io_device[14].port && io_device[14].id == DEV_NAME ? (3'b001 << io_device[14].num) : 3'b000) |
                      ((cpu_addr & io_device[15].mask) == io_device[15].port && io_device[15].id == DEV_NAME ? (3'b001 << io_device[15].num) : 3'b000);

endmodule
