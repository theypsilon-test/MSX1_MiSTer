module fdd #(parameter sysCLK, SECTORS=9, SECTOR_SIZE=512, TRACKS=80, TEST=0)
(
    input  logic            clk,
    input  logic            reset,
    FDD_if.FDD_mp           FDD_bus,

    //device config
    input logic       [3:0] speed,          // 0 - 300rpm / 1 - 360rpm
    input logic       [3:0] mfm,            // 0 - FM     / 1 - MFM
    //input logic       [3:0] sides,        // 0 - SS     / 1 - DS
    input logic       [1:0] density[4],     // 0 - 250kbit     / 1 - 500kbit    / 2 - 1000kbit
    input logic       [5:0] sectors[4],     // sectors per track
    input logic       [1:0] sector_size[4], // 0 - 128B / 1 - 256B / 2 - 512B / 3 - 1024B
    //hps image
    input logic       [3:0] img_mounted,
    input logic             img_readonly,
    input logic      [63:0] img_size,

    //SD block level access
    output logic     [31:0] sd_lba[0:3],
    output logic      [5:0] sd_blk_cnt[0:3],
    output logic      [3:0] sd_rd,
    output logic      [3:0] sd_wr,
    input  logic      [3:0] sd_ack,
   
    // SD byte level access. Signals for 2-PORT altsyncram.
    input  logic     [13:0] sd_buff_addr,
    input  logic      [7:0] sd_buff_dout,
    output logic      [7:0] sd_buff_din[0:3],
    input  logic            sd_buff_wr     
);

    
//https://map.grauw.nl/articles/low-level-disk/
//https://retrocmp.de/fdd/general/floppy-formats.htm

    logic motor_360rmp;
    clockEnabler #(.clkFreq(sysCLK), .targetFreq(6)) FDD_RPM360(
        .clk(clk),
        .en(motor_360rmp)
    );
    
    logic motor_300rmp;
    clockEnabler #(.clkFreq(sysCLK), .targetFreq(5)) FDD_RPM300(
        .clk(clk),
        .en(motor_300rmp)
    );

    logic msclk;
    clockEnabler #(.clkFreq(sysCLK), .targetFreq(1000)) FDD_MS(
        .clk(clk),
        .en(msclk)
    );

    logic bitRate_250;
    clockEnabler #(.clkFreq(sysCLK), .targetFreq(250000*2)) FDD_BITRATE_250(
        .clk(clk),
        .en(bitRate_250)
    );

    logic bitRate_500;
    clockEnabler #(.clkFreq(sysCLK), .targetFreq(500000*2)) FDD_BITRATE_500(
        .clk(clk),
        .en(bitRate_500)
    );

    logic bitRate_1000;
    clockEnabler #(.clkFreq(sysCLK), .targetFreq(1000000*2))  FDD_BITRATE_1000(
        .clk(clk),
        .en(bitRate_1000)
    );


    logic       drive_motor_rpm;
    logic       floppy_mfm;
    logic       floppy_sides;
    logic       floppy_bitRate;
    logic [5:0] floppy_sectors;
    logic [1:0] floppy_sectors_size;

    always_comb begin
        case (density[FDD_bus.USEL])
            2'd0: floppy_bitRate = bitRate_250;    
            2'd1: floppy_bitRate = bitRate_500;   
            2'd2: floppy_bitRate = bitRate_1000;
            default;
        endcase

        drive_motor_rpm     = speed[FDD_bus.USEL] ? motor_360rmp : motor_300rmp;
        floppy_mfm          = mfm[FDD_bus.USEL];
        floppy_sectors      = sectors[FDD_bus.USEL];
        floppy_sectors_size = sector_size[FDD_bus.USEL];
    end

    logic [3:0] motor_run;         // Stav motoru

    motor #(.TIMEOUTms(30000), .DELAYms(3)) FDD_motor(
        .clk(clk),
        .msclk(msclk),
        .reset(reset),
        .USEL(FDD_bus.USEL),
        .MOTORn(FDD_bus.MOTORn),
        .motor_run(motor_run)
    );

    //logic sides;
    ready FDD_ready(
        .clk(clk),
        .reset(reset),
        .USEL(FDD_bus.USEL),
        .motor_run(motor_run),
        .READYn(FDD_bus.READYn),
        .WPROTn(FDD_bus.WPROTn),
        .sides(/*sides*/),
        .img_mounted(img_mounted),
        .img_readonly(img_readonly),
        .img_size(img_size)
    );

    logic  [6:0] track;
    logic [12:0] buffer_addr;
    logic  [7:0] buffer_q;
    logic        track_ready;

    track #(.DELAYms(3), .MAX_TRACKS(80)) FDD_track(
        .clk(clk),
        .msclk(msclk),
        .reset(reset),
        .USEL(FDD_bus.USEL),
        .READYn(FDD_bus.READYn),
        .STEPn(FDD_bus.STEPn),
        .SDIRn(FDD_bus.SDIRn),
        .TRACK0n(FDD_bus.TRACK0n),
        .SIDEn(FDD_bus.SIDEn),
        
        .track(track),
        .disk_mounted(~FDD_bus.READYn),
        .disk_readonly(~FDD_bus.WPROTn),
        .disk_sides(/*sides*/),

        .track_ready(track_ready),
        .buffer_addr(buffer_addr),
        .buffer_q(buffer_q),

        .sd_lba(sd_lba),
        .sd_blk_cnt(sd_blk_cnt),
        .sd_rd(sd_rd),
        .sd_wr(sd_wr),
        .sd_ack(sd_ack),
        .sd_buff_addr(sd_buff_addr),
        .sd_buff_dout(sd_buff_dout),
        .sd_buff_din(sd_buff_din),
        .sd_buff_wr(sd_buff_wr)
    );

    transmit #(.sysCLK(sysCLK)) FDD_transmit(
        .clk(clk),
        .reset(reset),
        
        .drive_motor_rpm(drive_motor_rpm),
        .floppy_bitRate(floppy_bitRate),
        .floppy_mfm(floppy_mfm),
        .floppy_sectors(floppy_sectors),
        .floppy_sectors_size(floppy_sectors_size),

        //Track buffer
        .buffer_addr(buffer_addr),
        .buffer_q(buffer_q),
        .track_ready(track_ready),

        .track(track),
        .side(~FDD_bus.SIDEn),
        
        .INDEXn(FDD_bus.INDEXn),
        .READ_DATAn(FDD_bus.READ_DATAn)
    );

endmodule
